module mainn;
  initial 
    begin
      $display("Hello, World");
      $finish ;
    end
endmodule
