module axi4lite_read_fsm(clk, reset);

  //Input list
  input 	       clk, reset;

  //Output list

  //Signal declarations
  wire 	       clk, reset;

 //Add read/write state machine and connect up any other logic needed

endmodule // axi4lite_fsm
